-- Essas linhas devem estar em um arquivo  separado
-- File: meu_pkg.vhd
package meu_pkg is
  constant Nbit : natural := 2;
  type array1Dx1D is array (natural range <>) of bit_vector(Nbit-1 downto 0);
  type array2D is array (natural range <>, natural range <>) of bit;
end package;