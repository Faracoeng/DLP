-- FILE vector_adder.vhd --
---------------------------
configuration ifsc_cfg of vector_adder is
	-- for ifsc_v1 end for;
	for ifsc_v2 end for;
end configuration;